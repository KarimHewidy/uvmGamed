function void verify_test(GUVM_sequence_item cmd_trans,GUVM_result_transaction res_trans);
	
endfunction