`include "add.svh"